library verilog;
use verilog.vl_types.all;
entity lab6one_vlg_vec_tst is
end lab6one_vlg_vec_tst;
